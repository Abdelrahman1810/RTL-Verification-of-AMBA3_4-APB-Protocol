module APB_SVA();
    
endmodule